package wb_pkg;

endpackage
