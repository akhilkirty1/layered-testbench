// Specifies whether a transaction is a write or a read
typedef enum bit { READ, WRITE } i2c_op_t;
