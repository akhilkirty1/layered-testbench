mwglen@MattArch.4024