class i2cmb_env_configuration extends ncsu_env_configuration;

endclass
