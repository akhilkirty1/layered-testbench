// Determines whether a transaction is a write or a read
typedef enum bit { READ, WRITE } wb_op_t;
