class i2cmb_coverage extends ncsu_coverage;

endclass
