mwglen@MattArch.1806562331718805065