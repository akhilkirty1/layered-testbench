class wb_agent extends ncsu_agent;

endclass
