package i2c_pkg;
 typedef enum {READ, WRITE} i2c_op_t;
endpackage
