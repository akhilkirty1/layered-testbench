class wb_monitor extends ncsu_monitor;

endclass
