package i2cmb_env_pkg;
endpackage
