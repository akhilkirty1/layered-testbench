class wb_driver extends ncsu_driver;

endclass
