class i2cmb_generator extends ncsu_generator;

endclass
